module seven_seg_decoder(X0,X1,X2,X3,F);

	input X0, X1, X2, X3;
	output reg [0:6] F;
	
	always @(X0 or X1 or X2 or X3)
	begin
		case({X3, X2, X1, X0})
			4'b0000: F=7'b0000001;
			4'b0001: F=7'b1001111;
			4'b0010: F=7'b0010010;
			4'b0011: F=7'b0000110;
			4'b0100: F=7'b1001100;
			4'b0101: F=7'b0100100;
			4'b0110: F=7'b0100000;
			4'b0111: F=7'b0001111;
			4'b1000: F=7'b0000000;
			4'b1001: F=7'b0000100;
			4'b1010: F=7'b0001000;
			4'b1011: F=7'b1100000;
			4'b1100: F=7'b0110001;
			4'b1101: F=7'b1000010;
			4'b1110: F=7'b0110000;
			4'b1111: F=7'b0111000;
		endcase
	end
	
endmodule
